module main

import os { args }

fn main() {
	argument_parser := create_argument_parser(args[1..])
}